
//Verilog file of module adder


`timescale 1 ns / 1ns

module adder_net(operand_1,
operand_2,
NbarT, Si,
clk,
Sum, So);
input [0:31]operand_1;
input [0:31]operand_2;
input [0:0]clk;
output [0:31]Sum;
output So;
input NbarT;
input Si;

wire
adder_wire_1,
adder_wire_2,
adder_wire_3,
adder_wire_4,
adder_wire_5,
adder_wire_6,
adder_wire_7,
adder_wire_8,
adder_wire_9,
adder_wire_10,
adder_wire_11,
adder_wire_12,
adder_wire_13,
adder_wire_14,
adder_wire_15,
adder_wire_16,
adder_wire_17,
adder_wire_18,
adder_wire_19,
adder_wire_20,
adder_wire_21,
adder_wire_22,
adder_wire_23,
adder_wire_24,
adder_wire_25,
adder_wire_26,
adder_wire_27,
adder_wire_28,
adder_wire_29,
adder_wire_30,
adder_wire_31,
adder_wire_32,
adder_wire_33,
adder_wire_34,
adder_wire_35,
adder_wire_36,
adder_wire_37,
adder_wire_38,
adder_wire_39,
adder_wire_40,
adder_wire_41,
adder_wire_42,
adder_wire_43,
adder_wire_44,
adder_wire_45,
adder_wire_46,
adder_wire_47,
adder_wire_48,
adder_wire_49,
adder_wire_50,
adder_wire_51,
adder_wire_52,
adder_wire_53,
adder_wire_54,
adder_wire_55,
adder_wire_56,
adder_wire_57,
adder_wire_58,
adder_wire_59,
adder_wire_60,
adder_wire_61,
adder_wire_62,
adder_wire_63,
adder_wire_64,
adder_wire_65,
adder_wire_66,
adder_wire_67,
adder_wire_68,
adder_wire_69,
adder_wire_70,
adder_wire_71,
adder_wire_72,
adder_wire_73,
adder_wire_74,
adder_wire_75,
adder_wire_76,
adder_wire_77,
adder_wire_78,
adder_wire_79,
adder_wire_80,
adder_wire_81,
adder_wire_82,
adder_wire_83,
adder_wire_84,
adder_wire_85,
adder_wire_86,
adder_wire_87,
adder_wire_88,
adder_wire_89,
adder_wire_90,
adder_wire_91,
adder_wire_92,
adder_wire_93,
adder_wire_94,
adder_wire_95,
adder_wire_96,
adder_wire_97,
adder_wire_98,
adder_wire_99,
adder_wire_100,
adder_wire_101,
adder_wire_102,
adder_wire_103,
adder_wire_104,
adder_wire_105,
adder_wire_106,
adder_wire_107,
adder_wire_108,
adder_wire_109,
adder_wire_110,
adder_wire_111,
adder_wire_112,
adder_wire_113,
adder_wire_114,
adder_wire_115,
adder_wire_116,
adder_wire_117,
adder_wire_118,
adder_wire_119,
adder_wire_120,
adder_wire_121,
adder_wire_122,
adder_wire_123,
adder_wire_124,
adder_wire_125,
adder_wire_126,
adder_wire_127,
adder_wire_128,
adder_wire_129,
adder_wire_130,
adder_wire_131,
adder_wire_132,
adder_wire_133,
adder_wire_134,
adder_wire_135,
adder_wire_136,
adder_wire_137,
adder_wire_138,
adder_wire_139,
adder_wire_140,
adder_wire_141,
adder_wire_142,
adder_wire_143,
adder_wire_144,
adder_wire_145,
adder_wire_146,
adder_wire_147,
adder_wire_148,
adder_wire_149,
adder_wire_150,
adder_wire_151,
adder_wire_152,
adder_wire_153,
adder_wire_154,
adder_wire_155,
adder_wire_156,
adder_wire_157,
adder_wire_158,
adder_wire_159,
adder_wire_160,
adder_wire_161,
adder_wire_162,
adder_wire_163,
adder_wire_164,
adder_wire_165,
adder_wire_166,
adder_wire_167,
adder_wire_168,
adder_wire_169,
adder_wire_170,
adder_wire_171,
adder_wire_172,
adder_wire_173,
adder_wire_174,
adder_wire_175,
adder_wire_176,
adder_wire_177,
adder_wire_178,
adder_wire_179,
adder_wire_180,
adder_wire_181,
adder_wire_182,
adder_wire_183,
adder_wire_184,
adder_wire_185,
adder_wire_186,
adder_wire_187,
adder_wire_188,
adder_wire_189,
adder_wire_190,
adder_wire_191,
adder_wire_192,
adder_wire_193,
adder_wire_194,
adder_wire_195,
adder_wire_196,
adder_wire_197,
adder_wire_198,
adder_wire_199,
adder_wire_200,
adder_wire_201,
adder_wire_202,
adder_wire_203,
adder_wire_204,
adder_wire_205,
adder_wire_206,
adder_wire_207,
adder_wire_208,
adder_wire_209,
adder_wire_210,
adder_wire_211,
adder_wire_212,
adder_wire_213,
adder_wire_214,
adder_wire_215,
adder_wire_216,
adder_wire_217,
adder_wire_218,
adder_wire_219,
adder_wire_220,
adder_wire_221,
adder_wire_222,
adder_wire_223,
adder_wire_224,
adder_wire_225,
adder_wire_226,
adder_wire_227,
adder_wire_228,
adder_wire_229,
adder_wire_230,
adder_wire_231,
adder_wire_232,
adder_wire_233,
adder_wire_234,
adder_wire_235,
adder_wire_236,
adder_wire_237,
adder_wire_238,
adder_wire_239,
adder_wire_240,
adder_wire_241,
adder_wire_242,
adder_wire_243,
adder_wire_244,
adder_wire_245,
adder_wire_246,
adder_wire_247,
adder_wire_248,
adder_wire_249,
adder_wire_250,
adder_wire_251,
adder_wire_252,
adder_wire_253,
adder_wire_254,
adder_wire_255,
adder_wire_256,
adder_wire_257,
adder_wire_258,
adder_wire_259,
adder_wire_260,
adder_wire_261,
adder_wire_262,
adder_wire_263,
adder_wire_264,
adder_wire_265,
adder_wire_266,
adder_wire_267,
adder_wire_268,
adder_wire_269,
adder_wire_270,
adder_wire_271,
adder_wire_272,
adder_wire_273,
adder_wire_274,
adder_wire_275,
adder_wire_276,
adder_wire_277,
adder_wire_278,
adder_wire_279,
adder_wire_280,
adder_wire_281,
adder_wire_282,
adder_wire_283,
adder_wire_284,
adder_wire_285,
adder_wire_286,
adder_wire_287,
adder_wire_288,
adder_wire_289,
adder_wire_290,
adder_wire_291,
adder_wire_292,
adder_wire_293,
adder_wire_294,
adder_wire_29_0,
adder_wire_29_1,
adder_wire_26_0,
adder_wire_26_1,
adder_wire_32_0,
adder_wire_32_1,
adder_wire_35_0,
adder_wire_35_1,
adder_wire_38_0,
adder_wire_38_1,
adder_wire_68_0,
adder_wire_68_1,
adder_wire_68_2,
adder_wire_68_3,
adder_wire_68_4,
adder_wire_68_5,
adder_wire_68_6,
adder_wire_68_7,
adder_wire_68_8,
adder_wire_68_9,
adder_wire_68_10,
adder_wire_68_11,
adder_wire_68_12,
adder_wire_68_13,
adder_wire_68_14,
adder_wire_68_15,
adder_wire_68_16,
adder_wire_69_0,
adder_wire_69_1,
adder_wire_69_2,
adder_wire_69_3,
adder_wire_69_4,
adder_wire_69_5,
adder_wire_69_6,
adder_wire_69_7,
adder_wire_69_8,
adder_wire_69_9,
adder_wire_69_10,
adder_wire_69_11,
adder_wire_69_12,
adder_wire_69_13,
adder_wire_69_14,
adder_wire_69_15,
adder_wire_69_16,
adder_wire_20_0,
adder_wire_20_1,
adder_wire_20_2,
adder_wire_21_0,
adder_wire_21_1,
adder_wire_18_0,
adder_wire_18_1,
adder_wire_15_0,
adder_wire_15_1,
adder_wire_12_0,
adder_wire_12_1,
adder_wire_9_0,
adder_wire_9_1,
adder_wire_6_0,
adder_wire_6_1,
adder_wire_160_0,
adder_wire_160_1,
adder_wire_160_2,
adder_wire_160_3,
adder_wire_160_4,
adder_wire_160_5,
adder_wire_160_6,
adder_wire_160_7,
adder_wire_160_8,
adder_wire_160_9,
adder_wire_160_10,
adder_wire_160_11,
adder_wire_160_12,
adder_wire_160_13,
adder_wire_160_14,
adder_wire_160_15,
adder_wire_160_16,
adder_wire_160_17,
adder_wire_160_18,
adder_wire_160_19,
adder_wire_160_20,
adder_wire_160_21,
adder_wire_160_22,
adder_wire_204_0,
adder_wire_204_1,
adder_wire_204_2,
adder_wire_204_3,
adder_wire_204_4,
adder_wire_207_0,
adder_wire_207_1,
adder_wire_207_2,
adder_wire_207_3,
adder_wire_238_0,
adder_wire_238_1,
adder_wire_238_2,
adder_wire_238_3,
adder_wire_238_4,
adder_wire_238_5,
adder_wire_238_6,
adder_wire_238_7,
adder_wire_238_8,
adder_wire_238_9,
adder_wire_238_10,
adder_wire_238_11,
adder_wire_238_12,
adder_wire_238_13,
adder_wire_238_14,
adder_wire_238_15,
adder_wire_238_16,
adder_wire_241_0,
adder_wire_241_1,
adder_wire_241_2,
adder_wire_241_3,
adder_wire_241_4,
adder_wire_17_0,
adder_wire_17_1,
adder_wire_14_0,
adder_wire_14_1,
adder_wire_11_0,
adder_wire_11_1,
adder_wire_8_0,
adder_wire_8_1,
adder_wire_5_0,
adder_wire_5_1,
adder_wire_45_0,
adder_wire_45_1,
adder_wire_45_2,
adder_wire_45_3,
adder_wire_48_0,
adder_wire_48_1,
adder_wire_48_2,
adder_wire_48_3,
adder_wire_48_4,
adder_wire_48_5,
adder_wire_51_0,
adder_wire_51_1,
adder_wire_51_2,
adder_wire_51_3,
adder_wire_51_4,
adder_wire_51_5,
adder_wire_54_0,
adder_wire_54_1,
adder_wire_54_2,
adder_wire_54_3,
adder_wire_54_4,
adder_wire_54_5,
adder_wire_57_0,
adder_wire_57_1,
adder_wire_57_2,
adder_wire_57_3,
adder_wire_57_4,
adder_wire_57_5,
adder_wire_57_6,
adder_wire_57_7,
adder_wire_60_0,
adder_wire_60_1,
adder_wire_60_2,
adder_wire_60_3,
adder_wire_60_4,
adder_wire_60_5,
adder_wire_63_0,
adder_wire_63_1,
adder_wire_63_2,
adder_wire_63_3,
adder_wire_63_4,
adder_wire_63_5,
adder_wire_63_6,
adder_wire_63_7,
adder_wire_66_0,
adder_wire_66_1,
adder_wire_66_2,
adder_wire_66_3,
adder_wire_66_4,
adder_wire_66_5,
adder_wire_66_6,
adder_wire_66_7,
adder_wire_44_0,
adder_wire_44_1,
adder_wire_44_2,
adder_wire_44_3,
adder_wire_47_0,
adder_wire_47_1,
adder_wire_47_2,
adder_wire_47_3,
adder_wire_47_4,
adder_wire_47_5,
adder_wire_50_0,
adder_wire_50_1,
adder_wire_50_2,
adder_wire_50_3,
adder_wire_50_4,
adder_wire_50_5,
adder_wire_53_0,
adder_wire_53_1,
adder_wire_53_2,
adder_wire_53_3,
adder_wire_53_4,
adder_wire_53_5,
adder_wire_56_0,
adder_wire_56_1,
adder_wire_56_2,
adder_wire_56_3,
adder_wire_56_4,
adder_wire_56_5,
adder_wire_56_6,
adder_wire_56_7,
adder_wire_59_0,
adder_wire_59_1,
adder_wire_59_2,
adder_wire_59_3,
adder_wire_59_4,
adder_wire_59_5,
adder_wire_62_0,
adder_wire_62_1,
adder_wire_62_2,
adder_wire_62_3,
adder_wire_62_4,
adder_wire_62_5,
adder_wire_62_6,
adder_wire_62_7,
adder_wire_65_0,
adder_wire_65_1,
adder_wire_65_2,
adder_wire_65_3,
adder_wire_65_4,
adder_wire_65_5,
adder_wire_65_6,
adder_wire_65_7,
adder_wire_23_0,
adder_wire_23_1,
adder_wire_23_2,
adder_wire_24_0,
adder_wire_24_1,
adder_wire_27_0,
adder_wire_27_1,
adder_wire_30_0,
adder_wire_30_1,
adder_wire_33_0,
adder_wire_33_1,
adder_wire_36_0,
adder_wire_36_1,
adder_wire_39_0,
adder_wire_39_1;

pin #(65) pin_0 ({operand_1[0], operand_1[1], operand_1[2], operand_1[3], operand_1[4], operand_1[5], operand_1[6], operand_1[7], operand_1[8], operand_1[9], operand_1[10], operand_1[11], operand_1[12], operand_1[13], operand_1[14], operand_1[15], operand_1[16], operand_1[17], operand_1[18], operand_1[19], operand_1[20], operand_1[21], operand_1[22], operand_1[23], operand_1[24], operand_1[25], operand_1[26], operand_1[27], operand_1[28], operand_1[29], operand_1[30], operand_1[31], operand_2[0], operand_2[1], operand_2[2], operand_2[3], operand_2[4], operand_2[5], operand_2[6], operand_2[7], operand_2[8], operand_2[9], operand_2[10], operand_2[11], operand_2[12], operand_2[13], operand_2[14], operand_2[15], operand_2[16], operand_2[17], operand_2[18], operand_2[19], operand_2[20], operand_2[21], operand_2[22], operand_2[23], operand_2[24], operand_2[25], operand_2[26], operand_2[27], operand_2[28], operand_2[29], operand_2[30], operand_2[31], clk[0]}, {operand_1_0, operand_1_1, operand_1_2, operand_1_3, operand_1_4, operand_1_5, operand_1_6, operand_1_7, operand_1_8, operand_1_9, operand_1_10, operand_1_11, operand_1_12, operand_1_13, operand_1_14, operand_1_15, operand_1_16, operand_1_17, operand_1_18, operand_1_19, operand_1_20, operand_1_21, operand_1_22, operand_1_23, operand_1_24, operand_1_25, operand_1_26, operand_1_27, operand_1_28, operand_1_29, operand_1_30, operand_1_31, operand_2_0, operand_2_1, operand_2_2, operand_2_3, operand_2_4, operand_2_5, operand_2_6, operand_2_7, operand_2_8, operand_2_9, operand_2_10, operand_2_11, operand_2_12, operand_2_13, operand_2_14, operand_2_15, operand_2_16, operand_2_17, operand_2_18, operand_2_19, operand_2_20, operand_2_21, operand_2_22, operand_2_23, operand_2_24, operand_2_25, operand_2_26, operand_2_27, operand_2_28, operand_2_29, operand_2_30, operand_2_31, clk_0});

pout #(32) pout_0 ({Sum_0, Sum_1, Sum_2, Sum_3, Sum_4, Sum_5, Sum_6, Sum_7, Sum_8, Sum_9, Sum_10, Sum_11, Sum_12, Sum_13, Sum_14, Sum_15, Sum_16, Sum_17, Sum_18, Sum_19, Sum_20, Sum_21, Sum_22, Sum_23, Sum_24, Sum_25, Sum_26, Sum_27, Sum_28, Sum_29, Sum_30, Sum_31}, {Sum[0], Sum[1], Sum[2], Sum[3], Sum[4], Sum[5], Sum[6], Sum[7], Sum[8], Sum[9], Sum[10], Sum[11], Sum[12], Sum[13], Sum[14], Sum[15], Sum[16], Sum[17], Sum[18], Sum[19], Sum[20], Sum[21], Sum[22], Sum[23], Sum[24], Sum[25], Sum[26], Sum[27], Sum[28], Sum[29], Sum[30], Sum[31]});

fanout_n #(2, 0, 0) FANOUT_1 (adder_wire_29, {adder_wire_29_0, adder_wire_29_1});
fanout_n #(2, 0, 0) FANOUT_2 (adder_wire_26, {adder_wire_26_0, adder_wire_26_1});
fanout_n #(2, 0, 0) FANOUT_3 (adder_wire_32, {adder_wire_32_0, adder_wire_32_1});
fanout_n #(2, 0, 0) FANOUT_4 (adder_wire_35, {adder_wire_35_0, adder_wire_35_1});
fanout_n #(2, 0, 0) FANOUT_5 (adder_wire_38, {adder_wire_38_0, adder_wire_38_1});
fanout_n #(17, 0, 0) FANOUT_6 (adder_wire_68, {adder_wire_68_0, adder_wire_68_1, adder_wire_68_2, adder_wire_68_3, adder_wire_68_4, adder_wire_68_5, adder_wire_68_6, adder_wire_68_7, adder_wire_68_8, adder_wire_68_9, adder_wire_68_10, adder_wire_68_11, adder_wire_68_12, adder_wire_68_13, adder_wire_68_14, adder_wire_68_15, adder_wire_68_16});
fanout_n #(17, 0, 0) FANOUT_7 (adder_wire_69, {adder_wire_69_0, adder_wire_69_1, adder_wire_69_2, adder_wire_69_3, adder_wire_69_4, adder_wire_69_5, adder_wire_69_6, adder_wire_69_7, adder_wire_69_8, adder_wire_69_9, adder_wire_69_10, adder_wire_69_11, adder_wire_69_12, adder_wire_69_13, adder_wire_69_14, adder_wire_69_15, adder_wire_69_16});
fanout_n #(3, 0, 0) FANOUT_8 (adder_wire_20, {adder_wire_20_0, adder_wire_20_1, adder_wire_20_2});
fanout_n #(2, 0, 0) FANOUT_9 (adder_wire_21, {adder_wire_21_0, adder_wire_21_1});
fanout_n #(2, 0, 0) FANOUT_10 (adder_wire_18, {adder_wire_18_0, adder_wire_18_1});
fanout_n #(2, 0, 0) FANOUT_11 (adder_wire_15, {adder_wire_15_0, adder_wire_15_1});
fanout_n #(2, 0, 0) FANOUT_12 (adder_wire_12, {adder_wire_12_0, adder_wire_12_1});
fanout_n #(2, 0, 0) FANOUT_13 (adder_wire_9, {adder_wire_9_0, adder_wire_9_1});
fanout_n #(2, 0, 0) FANOUT_14 (adder_wire_6, {adder_wire_6_0, adder_wire_6_1});
fanout_n #(23, 0, 0) FANOUT_15 (adder_wire_160, {adder_wire_160_0, adder_wire_160_1, adder_wire_160_2, adder_wire_160_3, adder_wire_160_4, adder_wire_160_5, adder_wire_160_6, adder_wire_160_7, adder_wire_160_8, adder_wire_160_9, adder_wire_160_10, adder_wire_160_11, adder_wire_160_12, adder_wire_160_13, adder_wire_160_14, adder_wire_160_15, adder_wire_160_16, adder_wire_160_17, adder_wire_160_18, adder_wire_160_19, adder_wire_160_20, adder_wire_160_21, adder_wire_160_22});
fanout_n #(5, 0, 0) FANOUT_16 (adder_wire_204, {adder_wire_204_0, adder_wire_204_1, adder_wire_204_2, adder_wire_204_3, adder_wire_204_4});
fanout_n #(4, 0, 0) FANOUT_17 (adder_wire_207, {adder_wire_207_0, adder_wire_207_1, adder_wire_207_2, adder_wire_207_3});
fanout_n #(17, 0, 0) FANOUT_18 (adder_wire_238, {adder_wire_238_0, adder_wire_238_1, adder_wire_238_2, adder_wire_238_3, adder_wire_238_4, adder_wire_238_5, adder_wire_238_6, adder_wire_238_7, adder_wire_238_8, adder_wire_238_9, adder_wire_238_10, adder_wire_238_11, adder_wire_238_12, adder_wire_238_13, adder_wire_238_14, adder_wire_238_15, adder_wire_238_16});
fanout_n #(5, 0, 0) FANOUT_19 (adder_wire_241, {adder_wire_241_0, adder_wire_241_1, adder_wire_241_2, adder_wire_241_3, adder_wire_241_4});
fanout_n #(2, 0, 0) FANOUT_20 (adder_wire_17, {adder_wire_17_0, adder_wire_17_1});
fanout_n #(2, 0, 0) FANOUT_21 (adder_wire_14, {adder_wire_14_0, adder_wire_14_1});
fanout_n #(2, 0, 0) FANOUT_22 (adder_wire_11, {adder_wire_11_0, adder_wire_11_1});
fanout_n #(2, 0, 0) FANOUT_23 (adder_wire_8, {adder_wire_8_0, adder_wire_8_1});
fanout_n #(2, 0, 0) FANOUT_24 (adder_wire_5, {adder_wire_5_0, adder_wire_5_1});
fanout_n #(4, 0, 0) FANOUT_25 (adder_wire_45, {adder_wire_45_0, adder_wire_45_1, adder_wire_45_2, adder_wire_45_3});
fanout_n #(6, 0, 0) FANOUT_26 (adder_wire_48, {adder_wire_48_0, adder_wire_48_1, adder_wire_48_2, adder_wire_48_3, adder_wire_48_4, adder_wire_48_5});
fanout_n #(6, 0, 0) FANOUT_27 (adder_wire_51, {adder_wire_51_0, adder_wire_51_1, adder_wire_51_2, adder_wire_51_3, adder_wire_51_4, adder_wire_51_5});
fanout_n #(6, 0, 0) FANOUT_28 (adder_wire_54, {adder_wire_54_0, adder_wire_54_1, adder_wire_54_2, adder_wire_54_3, adder_wire_54_4, adder_wire_54_5});
fanout_n #(8, 0, 0) FANOUT_29 (adder_wire_57, {adder_wire_57_0, adder_wire_57_1, adder_wire_57_2, adder_wire_57_3, adder_wire_57_4, adder_wire_57_5, adder_wire_57_6, adder_wire_57_7});
fanout_n #(6, 0, 0) FANOUT_30 (adder_wire_60, {adder_wire_60_0, adder_wire_60_1, adder_wire_60_2, adder_wire_60_3, adder_wire_60_4, adder_wire_60_5});
fanout_n #(8, 0, 0) FANOUT_31 (adder_wire_63, {adder_wire_63_0, adder_wire_63_1, adder_wire_63_2, adder_wire_63_3, adder_wire_63_4, adder_wire_63_5, adder_wire_63_6, adder_wire_63_7});
fanout_n #(8, 0, 0) FANOUT_32 (adder_wire_66, {adder_wire_66_0, adder_wire_66_1, adder_wire_66_2, adder_wire_66_3, adder_wire_66_4, adder_wire_66_5, adder_wire_66_6, adder_wire_66_7});
fanout_n #(4, 0, 0) FANOUT_33 (adder_wire_44, {adder_wire_44_0, adder_wire_44_1, adder_wire_44_2, adder_wire_44_3});
fanout_n #(6, 0, 0) FANOUT_34 (adder_wire_47, {adder_wire_47_0, adder_wire_47_1, adder_wire_47_2, adder_wire_47_3, adder_wire_47_4, adder_wire_47_5});
fanout_n #(6, 0, 0) FANOUT_35 (adder_wire_50, {adder_wire_50_0, adder_wire_50_1, adder_wire_50_2, adder_wire_50_3, adder_wire_50_4, adder_wire_50_5});
fanout_n #(6, 0, 0) FANOUT_36 (adder_wire_53, {adder_wire_53_0, adder_wire_53_1, adder_wire_53_2, adder_wire_53_3, adder_wire_53_4, adder_wire_53_5});
fanout_n #(8, 0, 0) FANOUT_37 (adder_wire_56, {adder_wire_56_0, adder_wire_56_1, adder_wire_56_2, adder_wire_56_3, adder_wire_56_4, adder_wire_56_5, adder_wire_56_6, adder_wire_56_7});
fanout_n #(6, 0, 0) FANOUT_38 (adder_wire_59, {adder_wire_59_0, adder_wire_59_1, adder_wire_59_2, adder_wire_59_3, adder_wire_59_4, adder_wire_59_5});
fanout_n #(8, 0, 0) FANOUT_39 (adder_wire_62, {adder_wire_62_0, adder_wire_62_1, adder_wire_62_2, adder_wire_62_3, adder_wire_62_4, adder_wire_62_5, adder_wire_62_6, adder_wire_62_7});
fanout_n #(8, 0, 0) FANOUT_40 (adder_wire_65, {adder_wire_65_0, adder_wire_65_1, adder_wire_65_2, adder_wire_65_3, adder_wire_65_4, adder_wire_65_5, adder_wire_65_6, adder_wire_65_7});
fanout_n #(3, 0, 0) FANOUT_41 (adder_wire_23, {adder_wire_23_0, adder_wire_23_1, adder_wire_23_2});
fanout_n #(2, 0, 0) FANOUT_42 (adder_wire_24, {adder_wire_24_0, adder_wire_24_1});
fanout_n #(2, 0, 0) FANOUT_43 (adder_wire_27, {adder_wire_27_0, adder_wire_27_1});
fanout_n #(2, 0, 0) FANOUT_44 (adder_wire_30, {adder_wire_30_0, adder_wire_30_1});
fanout_n #(2, 0, 0) FANOUT_45 (adder_wire_33, {adder_wire_33_0, adder_wire_33_1});
fanout_n #(2, 0, 0) FANOUT_46 (adder_wire_36, {adder_wire_36_0, adder_wire_36_1});
fanout_n #(2, 0, 0) FANOUT_47 (adder_wire_39, {adder_wire_39_0, adder_wire_39_1});


xnor_n #(2, 0, 0) XNOR_1 (adder_wire_1, {adder_wire_2, adder_wire_3});
xnor_n #(2, 0, 0) XNOR_2 (adder_wire_4, {adder_wire_5_0, adder_wire_6_0});
xnor_n #(2, 0, 0) XNOR_3 (adder_wire_7, {adder_wire_8_0, adder_wire_9_0});
xnor_n #(2, 0, 0) XNOR_4 (adder_wire_10, {adder_wire_11_0, adder_wire_12_0});
xnor_n #(2, 0, 0) XNOR_5 (adder_wire_13, {adder_wire_14_0, adder_wire_15_0});
xnor_n #(2, 0, 0) XNOR_6 (adder_wire_16, {adder_wire_17_0, adder_wire_18_0});
xnor_n #(2, 0, 0) XNOR_7 (adder_wire_19, {adder_wire_20_0, adder_wire_21_0});
xor_n #(2, 0, 0) XOR_1 (adder_wire_22, {adder_wire_23_0, adder_wire_24_0});
xor_n #(2, 0, 0) XOR_2 (adder_wire_25, {adder_wire_26_0, adder_wire_27_0});
xor_n #(2, 0, 0) XOR_3 (adder_wire_28, {adder_wire_29_0, adder_wire_30_0});
xor_n #(2, 0, 0) XOR_4 (adder_wire_31, {adder_wire_32_0, adder_wire_33_0});
xor_n #(2, 0, 0) XOR_5 (adder_wire_34, {adder_wire_35_0, adder_wire_36_0});
xor_n #(2, 0, 0) XOR_6 (adder_wire_37, {adder_wire_38_0, adder_wire_39_0});
xor_n #(2, 0, 0) XOR_7 (adder_wire_40, {adder_wire_41, adder_wire_42});
xor_n #(2, 0, 0) XOR_8 (adder_wire_43, {adder_wire_44_0, adder_wire_45_0});
xor_n #(2, 0, 0) XOR_9 (adder_wire_46, {adder_wire_47_0, adder_wire_48_0});
xor_n #(2, 0, 0) XOR_10 (adder_wire_49, {adder_wire_50_0, adder_wire_51_0});
xor_n #(2, 0, 0) XOR_11 (adder_wire_52, {adder_wire_53_0, adder_wire_54_0});
xor_n #(2, 0, 0) XOR_12 (adder_wire_55, {adder_wire_56_0, adder_wire_57_0});
xor_n #(2, 0, 0) XOR_13 (adder_wire_58, {adder_wire_59_0, adder_wire_60_0});
xor_n #(2, 0, 0) XOR_14 (adder_wire_61, {adder_wire_62_0, adder_wire_63_0});
xor_n #(2, 0, 0) XOR_15 (adder_wire_64, {adder_wire_65_0, adder_wire_66_0});
and_n #(2, 0, 0) AND_1 (adder_wire_29, {adder_wire_26_1, adder_wire_27_1});
and_n #(2, 0, 0) AND_2 (adder_wire_26, {adder_wire_23_1, adder_wire_24_1});
and_n #(2, 0, 0) AND_3 (adder_wire_32, {adder_wire_29_1, adder_wire_30_1});
and_n #(2, 0, 0) AND_4 (adder_wire_35, {adder_wire_32_1, adder_wire_33_1});
and_n #(2, 0, 0) AND_5 (adder_wire_38, {adder_wire_35_1, adder_wire_36_1});
and_n #(2, 0, 0) AND_6 (adder_wire_41, {adder_wire_38_1, adder_wire_39_1});
or_n #(2, 0, 0) OR_1 (adder_wire_67, {adder_wire_68_0, adder_wire_69_0});
notg #(0, 0) NOT_1 (adder_wire_70, adder_wire_68_1);
or_n #(2, 0, 0) OR_2 (adder_wire_71, {adder_wire_68_2, adder_wire_69_1});
notg #(0, 0) NOT_2 (adder_wire_72, adder_wire_68_3);
or_n #(2, 0, 0) OR_3 (adder_wire_73, {adder_wire_68_4, adder_wire_69_2});
notg #(0, 0) NOT_3 (adder_wire_74, adder_wire_68_5);
or_n #(2, 0, 0) OR_4 (adder_wire_75, {adder_wire_68_6, adder_wire_69_3});
notg #(0, 0) NOT_4 (adder_wire_76, adder_wire_68_7);
or_n #(2, 0, 0) OR_5 (adder_wire_77, {adder_wire_68_8, adder_wire_69_4});
notg #(0, 0) NOT_5 (adder_wire_78, adder_wire_68_9);
or_n #(2, 0, 0) OR_6 (adder_wire_79, {adder_wire_68_10, adder_wire_69_5});
notg #(0, 0) NOT_6 (adder_wire_80, adder_wire_68_11);
or_n #(2, 0, 0) OR_7 (adder_wire_81, {adder_wire_68_12, adder_wire_69_6});
notg #(0, 0) NOT_7 (adder_wire_82, adder_wire_68_13);
or_n #(2, 0, 0) OR_8 (adder_wire_83, {adder_wire_68_14, adder_wire_69_7});
notg #(0, 0) NOT_8 (adder_wire_84, adder_wire_68_15);
nor_n #(8, 0, 0) NOR_1 (adder_wire_68, {adder_wire_58, adder_wire_55, adder_wire_64, adder_wire_49, adder_wire_46, adder_wire_43, adder_wire_52, adder_wire_61});
notg #(0, 0) NOT_9 (adder_wire_85, adder_wire_60_1);
and_n #(2, 0, 0) AND_7 (adder_wire_86, {adder_wire_85, adder_wire_59_1});
notg #(0, 0) NOT_10 (adder_wire_87, adder_wire_57_1);
and_n #(2, 0, 0) AND_8 (adder_wire_88, {adder_wire_87, adder_wire_56_1});
notg #(0, 0) NOT_11 (adder_wire_89, adder_wire_48_1);
and_n #(2, 0, 0) AND_9 (adder_wire_90, {adder_wire_89, adder_wire_47_1});
notg #(0, 0) NOT_12 (adder_wire_91, adder_wire_48_2);
or_n #(2, 0, 0) OR_9 (adder_wire_92, {adder_wire_91, adder_wire_47_2});
notg #(0, 0) NOT_13 (adder_wire_93, adder_wire_45_1);
and_n #(3, 0, 0) AND_10 (adder_wire_94, {adder_wire_93, adder_wire_92, adder_wire_44_1});
notg #(0, 0) NOT_14 (adder_wire_95, adder_wire_96);
and_n #(2, 0, 0) AND_11 (adder_wire_97, {adder_wire_95, adder_wire_98});
or_n #(4, 0, 0) OR_10 (adder_wire_99, {adder_wire_86, adder_wire_88, adder_wire_100, adder_wire_101});
and_n #(2, 0, 0) AND_12 (adder_wire_100, {adder_wire_102, adder_wire_62_1});
and_n #(2, 0, 0) AND_13 (adder_wire_101, {adder_wire_103, adder_wire_65_1});
or_n #(2, 0, 0) OR_11 (adder_wire_104, {adder_wire_105, adder_wire_56_2});
and_n #(3, 0, 0) AND_14 (adder_wire_106, {adder_wire_104, adder_wire_107, adder_wire_53_1});
or_n #(2, 0, 0) OR_12 (adder_wire_108, {adder_wire_109, adder_wire_53_2});
and_n #(2, 0, 0) AND_15 (adder_wire_110, {adder_wire_108, adder_wire_111});
notg #(0, 0) NOT_15 (adder_wire_102, adder_wire_63_1);
or_n #(2, 0, 0) OR_13 (adder_wire_111, {adder_wire_112, adder_wire_56_3});
and_n #(2, 0, 0) AND_16 (adder_wire_113, {adder_wire_114, adder_wire_50_1});
or_n #(2, 0, 0) OR_14 (adder_wire_115, {adder_wire_113, adder_wire_116});
or_n #(2, 0, 0) OR_15 (adder_wire_117, {adder_wire_118, adder_wire_50_2});
and_n #(2, 0, 0) AND_17 (adder_wire_116, {adder_wire_117, adder_wire_119});
or_n #(2, 0, 0) OR_16 (adder_wire_119, {adder_wire_90, adder_wire_94});
or_n #(2, 0, 0) OR_17 (adder_wire_98, {adder_wire_99, adder_wire_120});
or_n #(2, 0, 0) OR_18 (adder_wire_120, {adder_wire_106, adder_wire_121});
and_n #(2, 0, 0) AND_18 (adder_wire_121, {adder_wire_110, adder_wire_115});
notg #(0, 0) NOT_16 (adder_wire_103, adder_wire_66_1);
notg #(0, 0) NOT_17 (adder_wire_105, adder_wire_57_2);
notg #(0, 0) NOT_18 (adder_wire_107, adder_wire_54_1);
notg #(0, 0) NOT_19 (adder_wire_109, adder_wire_54_2);
notg #(0, 0) NOT_20 (adder_wire_112, adder_wire_57_3);
notg #(0, 0) NOT_21 (adder_wire_114, adder_wire_51_1);
notg #(0, 0) NOT_22 (adder_wire_118, adder_wire_51_2);
notg #(0, 0) NOT_23 (adder_wire_122, adder_wire_59_2);
and_n #(2, 0, 0) AND_19 (adder_wire_123, {adder_wire_122, adder_wire_60_2});
notg #(0, 0) NOT_24 (adder_wire_124, adder_wire_56_4);
and_n #(2, 0, 0) AND_20 (adder_wire_125, {adder_wire_124, adder_wire_57_4});
notg #(0, 0) NOT_25 (adder_wire_126, adder_wire_47_3);
and_n #(2, 0, 0) AND_21 (adder_wire_127, {adder_wire_126, adder_wire_48_3});
notg #(0, 0) NOT_26 (adder_wire_128, adder_wire_47_4);
or_n #(2, 0, 0) OR_19 (adder_wire_129, {adder_wire_128, adder_wire_48_4});
notg #(0, 0) NOT_27 (adder_wire_130, adder_wire_44_2);
and_n #(3, 0, 0) AND_22 (adder_wire_131, {adder_wire_130, adder_wire_129, adder_wire_45_2});
notg #(0, 0) NOT_28 (adder_wire_132, adder_wire_133);
and_n #(2, 0, 0) AND_23 (adder_wire_69, {adder_wire_132, adder_wire_134});
or_n #(4, 0, 0) OR_20 (adder_wire_135, {adder_wire_123, adder_wire_125, adder_wire_136, adder_wire_137});
and_n #(2, 0, 0) AND_24 (adder_wire_136, {adder_wire_138, adder_wire_63_2});
and_n #(2, 0, 0) AND_25 (adder_wire_137, {adder_wire_139, adder_wire_66_2});
or_n #(2, 0, 0) OR_21 (adder_wire_140, {adder_wire_141, adder_wire_57_5});
and_n #(3, 0, 0) AND_26 (adder_wire_142, {adder_wire_140, adder_wire_143, adder_wire_54_3});
or_n #(2, 0, 0) OR_22 (adder_wire_144, {adder_wire_145, adder_wire_54_4});
and_n #(2, 0, 0) AND_27 (adder_wire_146, {adder_wire_144, adder_wire_147});
notg #(0, 0) NOT_29 (adder_wire_138, adder_wire_62_2);
or_n #(2, 0, 0) OR_23 (adder_wire_147, {adder_wire_148, adder_wire_57_6});
and_n #(2, 0, 0) AND_28 (adder_wire_149, {adder_wire_150, adder_wire_51_3});
or_n #(2, 0, 0) OR_24 (adder_wire_151, {adder_wire_149, adder_wire_152});
or_n #(2, 0, 0) OR_25 (adder_wire_153, {adder_wire_154, adder_wire_51_4});
and_n #(2, 0, 0) AND_29 (adder_wire_152, {adder_wire_153, adder_wire_155});
or_n #(2, 0, 0) OR_26 (adder_wire_155, {adder_wire_127, adder_wire_131});
or_n #(2, 0, 0) OR_27 (adder_wire_134, {adder_wire_135, adder_wire_156});
or_n #(2, 0, 0) OR_28 (adder_wire_156, {adder_wire_142, adder_wire_157});
and_n #(2, 0, 0) AND_30 (adder_wire_157, {adder_wire_146, adder_wire_151});
notg #(0, 0) NOT_30 (adder_wire_139, adder_wire_65_2);
notg #(0, 0) NOT_31 (adder_wire_141, adder_wire_56_5);
notg #(0, 0) NOT_32 (adder_wire_143, adder_wire_53_3);
notg #(0, 0) NOT_33 (adder_wire_145, adder_wire_53_4);
notg #(0, 0) NOT_34 (adder_wire_148, adder_wire_56_6);
notg #(0, 0) NOT_35 (adder_wire_150, adder_wire_50_3);
notg #(0, 0) NOT_36 (adder_wire_154, adder_wire_50_4);
bufg #(0, 0) BUF_1 (adder_wire_158, 1'b1);
or_n #(2, 0, 0) OR_29 (adder_wire_133, {adder_wire_169, adder_wire_170});
notg #(0, 0) NOT_37 (adder_wire_171, adder_wire_66_3);
and_n #(2, 0, 0) AND_31 (adder_wire_170, {adder_wire_171, adder_wire_65_3});
and_n #(3, 0, 0) AND_32 (adder_wire_172, {adder_wire_173, adder_wire_174, adder_wire_59_3});
or_n #(2, 0, 0) OR_30 (adder_wire_175, {adder_wire_172, adder_wire_176});
and_n #(2, 0, 0) AND_33 (adder_wire_169, {adder_wire_175, adder_wire_177});
notg #(0, 0) NOT_38 (adder_wire_178, adder_wire_66_4);
or_n #(2, 0, 0) OR_31 (adder_wire_177, {adder_wire_178, adder_wire_65_4});
notg #(0, 0) NOT_39 (adder_wire_179, adder_wire_63_3);
and_n #(2, 0, 0) AND_34 (adder_wire_176, {adder_wire_179, adder_wire_62_3});
notg #(0, 0) NOT_40 (adder_wire_180, adder_wire_63_4);
or_n #(2, 0, 0) OR_32 (adder_wire_174, {adder_wire_180, adder_wire_62_4});
notg #(0, 0) NOT_41 (adder_wire_173, adder_wire_60_3);
or_n #(2, 0, 0) OR_33 (adder_wire_96, {adder_wire_181, adder_wire_182});
notg #(0, 0) NOT_42 (adder_wire_183, adder_wire_65_5);
and_n #(2, 0, 0) AND_35 (adder_wire_182, {adder_wire_183, adder_wire_66_5});
and_n #(3, 0, 0) AND_36 (adder_wire_184, {adder_wire_185, adder_wire_186, adder_wire_60_4});
or_n #(2, 0, 0) OR_34 (adder_wire_187, {adder_wire_184, adder_wire_188});
and_n #(2, 0, 0) AND_37 (adder_wire_181, {adder_wire_187, adder_wire_189});
notg #(0, 0) NOT_43 (adder_wire_190, adder_wire_65_6);
or_n #(2, 0, 0) OR_35 (adder_wire_189, {adder_wire_190, adder_wire_66_6});
notg #(0, 0) NOT_44 (adder_wire_191, adder_wire_62_5);
and_n #(2, 0, 0) AND_38 (adder_wire_188, {adder_wire_191, adder_wire_63_5});
notg #(0, 0) NOT_45 (adder_wire_192, adder_wire_62_6);
or_n #(2, 0, 0) OR_36 (adder_wire_186, {adder_wire_192, adder_wire_63_6});
notg #(0, 0) NOT_46 (adder_wire_185, adder_wire_59_4);
bufg #(0, 0) BUF_2 (Sum_31, adder_wire_160_0);
bufg #(0, 0) BUF_3 (Sum_21, adder_wire_160_1);
bufg #(0, 0) BUF_4 (Sum_20, adder_wire_160_2);
bufg #(0, 0) BUF_5 (Sum_19, adder_wire_160_3);
bufg #(0, 0) BUF_6 (Sum_18, adder_wire_160_4);
bufg #(0, 0) BUF_7 (Sum_17, adder_wire_160_5);
bufg #(0, 0) BUF_8 (Sum_16, adder_wire_160_6);
bufg #(0, 0) BUF_9 (Sum_15, adder_wire_160_7);
bufg #(0, 0) BUF_10 (Sum_14, adder_wire_160_8);
bufg #(0, 0) BUF_11 (Sum_13, adder_wire_160_9);
bufg #(0, 0) BUF_12 (Sum_12, adder_wire_160_10);
bufg #(0, 0) BUF_13 (Sum_30, adder_wire_160_11);
bufg #(0, 0) BUF_14 (Sum_11, adder_wire_160_12);
bufg #(0, 0) BUF_15 (Sum_10, adder_wire_160_13);
bufg #(0, 0) BUF_16 (Sum_9, adder_wire_160_14);
bufg #(0, 0) BUF_17 (Sum_8, adder_wire_193);
bufg #(0, 0) BUF_18 (Sum_7, adder_wire_194);
bufg #(0, 0) BUF_19 (Sum_6, adder_wire_195);
bufg #(0, 0) BUF_20 (Sum_5, adder_wire_196);
bufg #(0, 0) BUF_21 (Sum_4, adder_wire_197);
bufg #(0, 0) BUF_22 (Sum_3, adder_wire_198);
bufg #(0, 0) BUF_23 (Sum_2, adder_wire_199);
bufg #(0, 0) BUF_24 (Sum_29, adder_wire_160_15);
bufg #(0, 0) BUF_25 (Sum_1, adder_wire_200);
bufg #(0, 0) BUF_26 (Sum_0, adder_wire_201);
bufg #(0, 0) BUF_27 (Sum_28, adder_wire_160_16);
bufg #(0, 0) BUF_28 (Sum_27, adder_wire_160_17);
bufg #(0, 0) BUF_29 (Sum_26, adder_wire_160_18);
bufg #(0, 0) BUF_30 (Sum_25, adder_wire_160_19);
bufg #(0, 0) BUF_31 (Sum_24, adder_wire_160_20);
bufg #(0, 0) BUF_32 (Sum_23, adder_wire_160_21);
bufg #(0, 0) BUF_33 (Sum_22, adder_wire_160_22);
bufg #(0, 0) BUF_34 (adder_wire_160, 1'b0);
notg #(0, 0) NOT_47 (adder_wire_240, adder_wire_241_0);
and_n #(2, 0, 0) AND_39 (adder_wire_242, {adder_wire_241_1, adder_wire_204_0});
and_n #(3, 0, 0) AND_40 (adder_wire_235, {adder_wire_241_2, adder_wire_204_1, adder_wire_207_0});
and_n #(2, 0, 0) AND_41 (adder_wire_202, {adder_wire_241_3, adder_wire_243});
notg #(0, 0) NOT_48 (adder_wire_205, adder_wire_239);
nand_n #(2, 0, 0) NAND_1 (adder_wire_239, {adder_wire_204_2, adder_wire_241_4});
notg #(0, 0) NOT_49 (adder_wire_203, adder_wire_204_3);
nand_n #(2, 0, 0) NAND_2 (adder_wire_243, {adder_wire_204_4, adder_wire_207_1});
notg #(0, 0) NOT_50 (adder_wire_206, adder_wire_207_2);
notg #(0, 0) NOT_51 (adder_wire_244, adder_wire_207_3);
bufg #(0, 0) BUF_35 (adder_wire_159, clk_0);
or_n #(2, 0, 0) OR_37 (adder_wire_17, {adder_wire_20_1, adder_wire_21_1});
notg #(0, 0) NOT_52 (adder_wire_245, adder_wire_20_2);
or_n #(2, 0, 0) OR_38 (adder_wire_14, {adder_wire_18_1, adder_wire_17_1});
or_n #(2, 0, 0) OR_39 (adder_wire_11, {adder_wire_15_1, adder_wire_14_1});
or_n #(2, 0, 0) OR_40 (adder_wire_8, {adder_wire_12_1, adder_wire_11_1});
or_n #(2, 0, 0) OR_41 (adder_wire_5, {adder_wire_9_1, adder_wire_8_1});
or_n #(2, 0, 0) OR_42 (adder_wire_2, {adder_wire_6_1, adder_wire_5_1});
or_n #(2, 0, 0) OR_43 (adder_wire_161, {adder_wire_246, adder_wire_247});
and_n #(2, 0, 0) AND_42 (adder_wire_246, {adder_wire_245, adder_wire_238_0});
notg #(0, 0) NOT_53 (adder_wire_248, adder_wire_238_1);
and_n #(2, 0, 0) AND_43 (adder_wire_247, {adder_wire_248, adder_wire_224});
or_n #(2, 0, 0) OR_44 (adder_wire_162, {adder_wire_249, adder_wire_250});
and_n #(2, 0, 0) AND_44 (adder_wire_249, {adder_wire_19, adder_wire_238_2});
notg #(0, 0) NOT_54 (adder_wire_251, adder_wire_238_3);
and_n #(2, 0, 0) AND_45 (adder_wire_250, {adder_wire_251, adder_wire_222});
or_n #(2, 0, 0) OR_45 (adder_wire_163, {adder_wire_252, adder_wire_253});
and_n #(2, 0, 0) AND_46 (adder_wire_252, {adder_wire_16, adder_wire_238_4});
notg #(0, 0) NOT_55 (adder_wire_254, adder_wire_238_5);
and_n #(2, 0, 0) AND_47 (adder_wire_253, {adder_wire_254, adder_wire_220});
or_n #(2, 0, 0) OR_46 (adder_wire_164, {adder_wire_255, adder_wire_256});
and_n #(2, 0, 0) AND_48 (adder_wire_255, {adder_wire_13, adder_wire_238_6});
notg #(0, 0) NOT_56 (adder_wire_257, adder_wire_238_7);
and_n #(2, 0, 0) AND_49 (adder_wire_256, {adder_wire_257, adder_wire_218});
or_n #(2, 0, 0) OR_47 (adder_wire_165, {adder_wire_258, adder_wire_259});
and_n #(2, 0, 0) AND_50 (adder_wire_258, {adder_wire_10, adder_wire_238_8});
notg #(0, 0) NOT_57 (adder_wire_260, adder_wire_238_9);
and_n #(2, 0, 0) AND_51 (adder_wire_259, {adder_wire_260, adder_wire_216});
or_n #(2, 0, 0) OR_48 (adder_wire_166, {adder_wire_261, adder_wire_262});
and_n #(2, 0, 0) AND_52 (adder_wire_261, {adder_wire_7, adder_wire_238_10});
notg #(0, 0) NOT_58 (adder_wire_263, adder_wire_238_11);
and_n #(2, 0, 0) AND_53 (adder_wire_262, {adder_wire_263, adder_wire_214});
or_n #(2, 0, 0) OR_49 (adder_wire_167, {adder_wire_264, adder_wire_265});
and_n #(2, 0, 0) AND_54 (adder_wire_264, {adder_wire_4, adder_wire_238_12});
notg #(0, 0) NOT_59 (adder_wire_266, adder_wire_238_13);
and_n #(2, 0, 0) AND_55 (adder_wire_265, {adder_wire_266, adder_wire_212});
or_n #(2, 0, 0) OR_50 (adder_wire_168, {adder_wire_267, adder_wire_268});
and_n #(2, 0, 0) AND_56 (adder_wire_267, {adder_wire_1, adder_wire_238_14});
notg #(0, 0) NOT_60 (adder_wire_269, adder_wire_238_15);
and_n #(2, 0, 0) AND_57 (adder_wire_268, {adder_wire_269, adder_wire_210});
and_n #(2, 0, 0) AND_58 (adder_wire_208, {adder_wire_242, adder_wire_244});
bufg #(0, 0) BUF_36 (adder_wire_45, operand_1_8);
bufg #(0, 0) BUF_37 (adder_wire_48, operand_1_7);
bufg #(0, 0) BUF_38 (adder_wire_51, operand_1_6);
bufg #(0, 0) BUF_39 (adder_wire_54, operand_1_5);
bufg #(0, 0) BUF_40 (adder_wire_57, operand_1_4);
bufg #(0, 0) BUF_41 (adder_wire_60, operand_1_3);
bufg #(0, 0) BUF_42 (adder_wire_63, operand_1_2);
bufg #(0, 0) BUF_43 (adder_wire_66, operand_1_1);
bufg #(0, 0) BUF_44 (adder_wire_236, operand_1_0);
and_n #(2, 0, 0) AND_59 (adder_wire_270, {adder_wire_45_3, adder_wire_83});
and_n #(2, 0, 0) AND_60 (adder_wire_271, {adder_wire_48_5, adder_wire_81});
and_n #(2, 0, 0) AND_61 (adder_wire_272, {adder_wire_51_5, adder_wire_79});
and_n #(2, 0, 0) AND_62 (adder_wire_273, {adder_wire_54_5, adder_wire_77});
and_n #(2, 0, 0) AND_63 (adder_wire_274, {adder_wire_57_7, adder_wire_75});
and_n #(2, 0, 0) AND_64 (adder_wire_275, {adder_wire_60_5, adder_wire_73});
and_n #(2, 0, 0) AND_65 (adder_wire_276, {adder_wire_63_7, adder_wire_71});
and_n #(2, 0, 0) AND_66 (adder_wire_277, {adder_wire_66_7, adder_wire_67});
bufg #(0, 0) BUF_45 (adder_wire_44, operand_2_8);
bufg #(0, 0) BUF_46 (adder_wire_47, operand_2_7);
bufg #(0, 0) BUF_47 (adder_wire_50, operand_2_6);
bufg #(0, 0) BUF_48 (adder_wire_53, operand_2_5);
bufg #(0, 0) BUF_49 (adder_wire_56, operand_2_4);
bufg #(0, 0) BUF_50 (adder_wire_59, operand_2_3);
bufg #(0, 0) BUF_51 (adder_wire_62, operand_2_2);
bufg #(0, 0) BUF_52 (adder_wire_65, operand_2_1);
and_n #(3, 0, 0) AND_67 (adder_wire_278, {adder_wire_44_3, adder_wire_84, adder_wire_279});
and_n #(3, 0, 0) AND_68 (adder_wire_280, {adder_wire_47_5, adder_wire_82, adder_wire_281});
and_n #(3, 0, 0) AND_69 (adder_wire_282, {adder_wire_50_5, adder_wire_80, adder_wire_283});
and_n #(3, 0, 0) AND_70 (adder_wire_284, {adder_wire_53_5, adder_wire_78, adder_wire_285});
and_n #(3, 0, 0) AND_71 (adder_wire_286, {adder_wire_56_7, adder_wire_76, adder_wire_287});
and_n #(3, 0, 0) AND_72 (adder_wire_288, {adder_wire_59_5, adder_wire_74, adder_wire_289});
and_n #(3, 0, 0) AND_73 (adder_wire_290, {adder_wire_62_7, adder_wire_72, adder_wire_291});
and_n #(3, 0, 0) AND_74 (adder_wire_292, {adder_wire_65_7, adder_wire_70, adder_wire_293});
notg #(0, 0) NOT_61 (adder_wire_237, adder_wire_238_16);
notg #(0, 0) NOT_62 (adder_wire_225, adder_wire_294);
nor_n #(3, 0, 0) NOR_2 (adder_wire_294, {adder_wire_69_8, adder_wire_97, adder_wire_68_16});
notg #(0, 0) NOT_63 (adder_wire_293, adder_wire_69_9);
notg #(0, 0) NOT_64 (adder_wire_291, adder_wire_69_10);
notg #(0, 0) NOT_65 (adder_wire_289, adder_wire_69_11);
notg #(0, 0) NOT_66 (adder_wire_287, adder_wire_69_12);
notg #(0, 0) NOT_67 (adder_wire_285, adder_wire_69_13);
notg #(0, 0) NOT_68 (adder_wire_283, adder_wire_69_14);
notg #(0, 0) NOT_69 (adder_wire_281, adder_wire_69_15);
notg #(0, 0) NOT_70 (adder_wire_279, adder_wire_69_16);
notg #(0, 0) NOT_71 (adder_wire_233, adder_wire_23_2);
or_n #(2, 0, 0) OR_51 (adder_wire_23, {adder_wire_270, adder_wire_278});
or_n #(2, 0, 0) OR_52 (adder_wire_24, {adder_wire_271, adder_wire_280});
or_n #(2, 0, 0) OR_53 (adder_wire_27, {adder_wire_272, adder_wire_282});
or_n #(2, 0, 0) OR_54 (adder_wire_30, {adder_wire_273, adder_wire_284});
or_n #(2, 0, 0) OR_55 (adder_wire_33, {adder_wire_274, adder_wire_286});
or_n #(2, 0, 0) OR_56 (adder_wire_36, {adder_wire_275, adder_wire_288});
or_n #(2, 0, 0) OR_57 (adder_wire_39, {adder_wire_276, adder_wire_290});
or_n #(2, 0, 0) OR_58 (adder_wire_42, {adder_wire_277, adder_wire_292});
dff DFF_1  (adder_wire_20, adder_wire_161, adder_wire_159, adder_wire_160, 1'b0, adder_wire_158, NbarT,Si, 1'b0);
dff DFF_2  (adder_wire_21, adder_wire_162, adder_wire_159, adder_wire_160, 1'b0, adder_wire_158, NbarT,adder_wire_20, 1'b0);
dff DFF_3  (adder_wire_18, adder_wire_163, adder_wire_159, adder_wire_160, 1'b0, adder_wire_158, NbarT,adder_wire_21, 1'b0);
dff DFF_4  (adder_wire_15, adder_wire_164, adder_wire_159, adder_wire_160, 1'b0, adder_wire_158, NbarT,adder_wire_18, 1'b0);
dff DFF_5  (adder_wire_12, adder_wire_165, adder_wire_159, adder_wire_160, 1'b0, adder_wire_158, NbarT,adder_wire_15, 1'b0);
dff DFF_6  (adder_wire_9, adder_wire_166, adder_wire_159, adder_wire_160, 1'b0, adder_wire_158, NbarT,adder_wire_12,  1'b0);
dff DFF_7  (adder_wire_6, adder_wire_167, adder_wire_159, adder_wire_160, 1'b0, adder_wire_158, NbarT,adder_wire_9,  1'b0);
dff DFF_8  (adder_wire_3, adder_wire_168, adder_wire_159, adder_wire_160, 1'b0, adder_wire_158, NbarT,adder_wire_6,  1'b0);
dff DFF_9  (adder_wire_204, adder_wire_203, adder_wire_159, adder_wire_160, 1'b0, adder_wire_202, NbarT,adder_wire_3,  1'b0);
dff DFF_10  (adder_wire_207, adder_wire_206, adder_wire_159, adder_wire_160, 1'b0, adder_wire_205, NbarT,adder_wire_204, 1'b0);
dff DFF_11  (adder_wire_210, adder_wire_209, adder_wire_159, adder_wire_160, 1'b0, adder_wire_208, NbarT,adder_wire_207, 1'b0);
dff DFF_12  (adder_wire_212, adder_wire_211, adder_wire_159, adder_wire_160, 1'b0, adder_wire_208, NbarT,adder_wire_210, 1'b0);
dff DFF_13  (adder_wire_214, adder_wire_213, adder_wire_159, adder_wire_160, 1'b0, adder_wire_208, NbarT,adder_wire_212, 1'b0);
dff DFF_14  (adder_wire_216, adder_wire_215, adder_wire_159, adder_wire_160, 1'b0, adder_wire_208, NbarT,adder_wire_214, 1'b0);
dff DFF_15  (adder_wire_218, adder_wire_217, adder_wire_159, adder_wire_160, 1'b0, adder_wire_208, NbarT,adder_wire_216, 1'b0);
dff DFF_16  (adder_wire_220, adder_wire_219, adder_wire_159, adder_wire_160, 1'b0, adder_wire_208, NbarT,adder_wire_218, 1'b0);
dff DFF_17  (adder_wire_222, adder_wire_221, adder_wire_159, adder_wire_160, 1'b0, adder_wire_208, NbarT,adder_wire_220, 1'b0);
dff DFF_18  (adder_wire_224, adder_wire_223, adder_wire_159, adder_wire_160, 1'b0, adder_wire_208, NbarT,adder_wire_222, 1'b0);
dff DFF_19  (adder_wire_226, adder_wire_40, adder_wire_159, adder_wire_160, 1'b0, adder_wire_225, NbarT,adder_wire_224,  1'b0);
dff DFF_20  (adder_wire_227, adder_wire_37, adder_wire_159, adder_wire_160, 1'b0, adder_wire_225, NbarT,adder_wire_226,  1'b0);
dff DFF_21  (adder_wire_228, adder_wire_34, adder_wire_159, adder_wire_160, 1'b0, adder_wire_225, NbarT,adder_wire_227,  1'b0);
dff DFF_22  (adder_wire_229, adder_wire_31, adder_wire_159, adder_wire_160, 1'b0, adder_wire_225, NbarT,adder_wire_228,  1'b0);
dff DFF_23  (adder_wire_230, adder_wire_28, adder_wire_159, adder_wire_160, 1'b0, adder_wire_225, NbarT,adder_wire_229,  1'b0);
dff DFF_24  (adder_wire_231, adder_wire_25, adder_wire_159, adder_wire_160, 1'b0, adder_wire_225, NbarT,adder_wire_230,  1'b0);
dff DFF_25  (adder_wire_232, adder_wire_22, adder_wire_159, adder_wire_160, 1'b0, adder_wire_225, NbarT,adder_wire_231,  1'b0);
dff DFF_26  (adder_wire_234, adder_wire_233, adder_wire_159, adder_wire_160, 1'b0, adder_wire_225, NbarT,adder_wire_232, 1'b0);
dff DFF_27  (adder_wire_201, adder_wire_236, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_234, 1'b0);
dff DFF_28  (adder_wire_200, adder_wire_3, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_201,  1'b0);
dff DFF_29  (adder_wire_199, adder_wire_6, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_200,  1'b0);
dff DFF_30  (adder_wire_198, adder_wire_9, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_199,  1'b0);
dff DFF_31  (adder_wire_197, adder_wire_12, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_198,  1'b0);
dff DFF_32  (adder_wire_196, adder_wire_15, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_197,  1'b0);
dff DFF_33  (adder_wire_195, adder_wire_18, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_196,  1'b0);
dff DFF_34  (adder_wire_194, adder_wire_21, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_195,  1'b0);
dff DFF_35  (adder_wire_193, adder_wire_20, adder_wire_159, adder_wire_160, 1'b0, adder_wire_235, NbarT,adder_wire_194,  1'b0);
dff DFF_36  (adder_wire_238, adder_wire_237, adder_wire_159, adder_wire_160, 1'b0, adder_wire_237, NbarT,adder_wire_193, 1'b0);
dff DFF_37  (adder_wire_241, adder_wire_240, adder_wire_159, adder_wire_160, 1'b0, adder_wire_239, NbarT,adder_wire_238, 1'b0);
dff DFF_38  (adder_wire_223, adder_wire_234, adder_wire_159, 1'b0, 1'b0, 1'b1, NbarT,adder_wire_241, 1'b0);
dff DFF_39  (adder_wire_221, adder_wire_232, adder_wire_159, 1'b0, 1'b0, 1'b1, NbarT,adder_wire_223, 1'b0);
dff DFF_40  (adder_wire_219, adder_wire_231, adder_wire_159, 1'b0, 1'b0, 1'b1, NbarT,adder_wire_221, 1'b0);
dff DFF_41  (adder_wire_217, adder_wire_230, adder_wire_159, 1'b0, 1'b0, 1'b1, NbarT,adder_wire_219, 1'b0);
dff DFF_42  (adder_wire_215, adder_wire_229, adder_wire_159, 1'b0, 1'b0, 1'b1, NbarT,adder_wire_217, 1'b0);
dff DFF_43  (adder_wire_213, adder_wire_228, adder_wire_159, 1'b0, 1'b0, 1'b1, NbarT,adder_wire_215, 1'b0);
dff DFF_44  (adder_wire_211, adder_wire_227, adder_wire_159, 1'b0, 1'b0, 1'b1, NbarT,adder_wire_213, 1'b0);
dff DFF_45  (adder_wire_209, adder_wire_226, adder_wire_159, 1'b0, 1'b0, 1'b1, NbarT,adder_wire_211, 1'b0);

assign So = adder_wire_209;
endmodule
